// pseudocode of hft algorithm
